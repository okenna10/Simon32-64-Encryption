//NumStages defines the number of pipeline stages in Your design. Minimum Numstags = 1 is for non-pipelined design 
//i.e. no intermediate flip-flops between I/O flipflops.
localparam NumStages = 1;
// clock period in ns (nano second)
localparam ClkPeriod = 2;

